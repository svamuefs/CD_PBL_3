module comparator (
    
);
    
endmodule