module automacao (
	input a ,
	output b

);

endmodule